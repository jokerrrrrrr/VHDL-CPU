----------------------------------------------------------------------------------
-- Digitalteknik portef�lje 2
-- VHDL-CPU
-- Af Kent Stark Olsen og Leon Bonde Larsen
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity cpu is port 
		(
			clock: in std_logic
		); 
end cpu;

--architecture cpu_core of cpu is


--end cpu_core;